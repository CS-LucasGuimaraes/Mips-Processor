`timescale 1ps/1ps

module ctrl_unit (
    input [31:0] instr
);

