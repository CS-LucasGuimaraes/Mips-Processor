//////////////////////////
////// Instruções R //////
//////////////////////////

`define R_TYPE  6'b000000

`define JUMP    6'b00100X
`define JR      6'b001000

//////////////////////////
////// Instruções I //////
//////////////////////////

`define ADDI    6'b001000
`define BNE     6'b000101
`define LW      6'b100011
`define SW      6'b101011

//////////////////////////   
////// Instruções J //////
//////////////////////////

`define JAL     6'b000011